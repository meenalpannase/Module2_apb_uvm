`ifdef SEQUENCER
`define SEQUENCER
//include files 

//Import the UVM package
//class declaration

`endif
