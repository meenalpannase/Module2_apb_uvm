`ifdef DRV
`define DRV
//include files

//Importing the UVM package

class m_driver extends uvm_driver #(m_seq_item);
   //Declaring the virtual interface
  
   //Constructor
   
   
   //Build phase
  

   //Run phase
   
endclass
`endif
