`ifdef SEQ_ITEM
`define SEQ_ITEM
//Adding the UVM macros

//Importing the UVM package

class m_seq_item extends uvm_sequence_item;
   //variable declaration
   
   //Utility macros
  

   //Constructor
   
endclass
`endif
