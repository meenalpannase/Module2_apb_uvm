interface intf(input bit pclk,input bit prst);
   

   //Cloking block for driver
   
      //Default input and output declaration
      
   endclocking

   //Clocking block for monitor
  
      //Default input and output declaration
      
   endclocking

   //Modport declarations
  
endinterface

