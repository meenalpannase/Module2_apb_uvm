`ifdef 
`define
package test_pkg;
   //include and import uvm_macros ,pkg and files
  
endpackage
`endif
