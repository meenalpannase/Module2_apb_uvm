`ifdef TEST
`define TEST
//include files
"
//Importing the UVM package

class apb_test extends uvm_test;
  
   //s_sequence sseq;

   //Constructor
   

   //Build phase
   
 

   //Connect phase
  

   //Run phase
   

   //Write test case
  

   //Read test case
  
endclass
`endif
