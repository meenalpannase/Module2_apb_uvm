`ifdef MASTER_PACKAGE
`define MASTER_PACKAGE
package master_pkg;
   `include "uvm_macros.svh"
   import uvm_pkg::*;
  //include master files
endpackage
`endif
