`define addrWidth 
`define dataWidth 
