`ifdef SCOREBOARD
`define SCOREBOARD
//include files 


//Importing the UVM package

class apb_scoreboard extends uvm_scoreboard;


   //decalre analysis ports 

   //Constructor


   //Build phase
  

   //Connect Phase


   //Writing the data from driver
 

   //Writing the data from monitor
 

   //Run phase


   //Check phase
  

   //Report phase
 
endclass
`endif

