`ifdef AGENTM
`define AGENTM
//include files

class m_agent extends uvm_agent;
  
   //UVM Macros
  
   
   //constructor
   

   //Build Phase
   
   //Connect Phase
   
endclass
`endif
