`ifdef ENVIRONMENT
`define ENVIRONMENT
//include files

//Importing the UVM package

class apb_environment extends uvm_env;
  

   //Virtual Interface
 

  

   //Build phase
   

   //Connect phase
   
   //Run phase
  
endclass
`endif
