//define timescale

//include all files

//Importing UVM package

module apb_tbtop(); 
   //Clock and reset signal declaration
   
   //Interface instance
   
   //Clock generation
  
   //reset generation
   
   //DUT instance
  //set virtual interface
   
   initial 
   begin
      $dumpfile("dump.vcd"); 
      $dumpvars;
   end
endmodule
